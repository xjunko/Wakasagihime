module object

pub struct Spinner {
	HitObject
}
