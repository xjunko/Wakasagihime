module main

// vfmt off
import beatmap
// vfmt on

fn main() {
	beatmap.parse('/run/media/junko/2nd/Projects/Echidna/src/wakasagihime/sekai/assets/maps/poemdoll/master.sus')
}
