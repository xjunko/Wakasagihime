module objects

import wakasagihime.diva.beatmap.opcodes

pub struct BaseNode {
pub mut:
	commands opcodes.OPCode
}
